module testIf(clk,A,B);
input clk;
output reg [3:0] A+4'h0;
output reg [3:0] B=4'h0;
module testIf(clk,A,B);

module testIf(clk,A,B);
input clk;
output reg [3:0] A+4'h0;
output reg [3:0] B=4'h0;
