module test(x);
//test
//
//
//
//
endmodule
